`timescale 1ns / 1ns
module tb_top;

reg clk;
reg rst;

reg [7:0] mem[65535:0];
integer i;
integer f;

initial forever #5 clk = ~clk;

initial
begin
    $vcdplusfile("wave.vpd");
    $vcdpluson();
end

initial
begin
    // Reset
    clk = 0;
    rst = 1;
    repeat (5) @(posedge clk);
    rst = 0;

    // Load TCM memory
    for (i=0;i<65535;i=i+1)
        mem[i] = 0;

    f = $fopen("./app_test/app_test.bin", "r");
    i = $fread(mem, f);
    for (i=0;i<65535;i=i+1)
        u_mem.write(i, mem[i]);
    
    repeat(30000) @(posedge clk);
    $finish;
end

wire          mem_i_rd_w;
wire [ 31:0]  mem_i_pc_w;
wire [ 31:0]  mem_d_addr_w;
wire [ 31:0]  mem_d_data_wr_w;
wire          mem_d_rd_w;
wire [  3:0]  mem_d_wr_w;
wire          mem_i_accept_w;
wire          mem_i_valid_w;
wire [ 31:0]  mem_i_inst_w;
wire [ 31:0]  mem_d_data_rd_w;
wire          mem_d_accept_w;
wire          mem_d_ack_w;

uriscv_core u_dut (
    .clk_i(clk),
    .rst_i(rst),
    .mem_d_data_rd_i(mem_d_data_rd_w),
    .mem_d_accept_i(mem_d_accept_w),
    .mem_d_ack_i(mem_d_ack_w),
    .mem_i_accept_i(mem_i_accept_w),
    .mem_i_valid_i(mem_i_valid_w),
    .mem_i_inst_i(mem_i_inst_w),
    .intr_i(1'b0),
    .reset_vector_i(32'h0),
    .cpu_id_i('b0),
    .mem_d_addr_o(mem_d_addr_w),
    .mem_d_data_wr_o(mem_d_data_wr_w),
    .mem_d_rd_o(mem_d_rd_w),
    .mem_d_wr_o(mem_d_wr_w),
    .mem_i_rd_o(mem_i_rd_w),
    .mem_i_pc_o(mem_i_pc_w)
);

tcm_mem u_mem (
    .clk_i(clk),
    .rst_i(rst),
    .mem_i_rd_i(mem_i_rd_w),
    .mem_i_flush_i(1'b0),
    .mem_i_invalidate_i(1'b0),
    .mem_i_pc_i(mem_i_pc_w),
    .mem_d_addr_i(mem_d_addr_w),
    .mem_d_data_wr_i(mem_d_data_wr_w),
    .mem_d_rd_i(mem_d_rd_w),
    .mem_d_wr_i(mem_d_wr_w),
    .mem_d_cacheable_i(1'b0),
    .mem_d_req_tag_i(11'h0),
    .mem_d_invalidate_i(1'b0),
    .mem_d_writeback_i(1'b0),
    .mem_d_flush_i(1'b0),
    .mem_i_accept_o(mem_i_accept_w),
    .mem_i_valid_o(mem_i_valid_w),
    .mem_i_error_o(),
    .mem_i_inst_o(mem_i_inst_w),
    .mem_d_data_rd_o(mem_d_data_rd_w),
    .mem_d_accept_o(mem_d_accept_w),
    .mem_d_ack_o(mem_d_ack_w),
    .mem_d_error_o(),
    .mem_d_resp_tag_o()
);

endmodule
